module nor_gate_st(
    input a,
    input b,
    output y
);

nor(y,a,b);

endmodule