module xor_gate_st(
    input a,
    input b,
    output y
);

xor(y,a,b);

endmodule