module or_gate_st(
    input a,
    input b,
    output y
);

or(y,a,b);

endmodule

