module nand_gate_st(
    input a,
    input b,
    output y
);

nand(y,a,b);

endmodule