module and_gate_st(
    input a,
    input b,
    output y
);

and(y,a,b);

endmodule
