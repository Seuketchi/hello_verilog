module xnor_gate_st(
    input a,
    input b,
    output y
);

xnor(y,a,b);

endmodule