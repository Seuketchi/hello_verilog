module not_gate_st(
    input a,
    output y
);

not(y,a);

endmodule