module not_gate_df(
    input a,
    output y
);
    assign y = ~a;
endmodule