module seven_segment_display(
    input [15:0] i,
    output reg [6:0] y
);

always @(*) begin
    case (i)
            16'b0000_0000_0000_0001: y = 7'b0111111; // 0
            16'b0000_0000_0000_0010: y = 7'b0000110; // 1
            16'b0000_0000_0000_0100: y = 7'b1011011; // 2
            16'b0000_0000_0000_1000: y = 7'b1001111; // 3
            16'b0000_0000_0001_0000: y = 7'b1100110; // 4
            16'b0000_0000_0010_0000: y = 7'b1101101; // 5
            16'b0000_0000_0100_0000: y = 7'b1111101; // 6
            16'b0000_0000_1000_0000: y = 7'b0000111; // 7
            16'b0000_0001_0000_0000: y = 7'b1111111; // 8
            16'b0000_0010_0000_0000: y = 7'b1101111; // 9
            16'b0000_0100_0000_0000: y = 7'b1110111; // A
            16'b0000_1000_0000_0000: y = 7'b1111100; // B
            16'b0001_0000_0000_0000: y = 7'b0111001; // C
            16'b0010_0000_0000_0000: y = 7'b1011110; // D
            16'b0100_0000_0000_0000: y = 7'b1111001; // E
            16'b1000_0000_0000_0000: y = 7'b1110001; // F
            default: y = 7'b0000000; // Off
    endcase
end

endmodule